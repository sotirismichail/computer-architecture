library IEEE;
use IEEE.STD_LOGIC_1164.all;

package array_5bit is
	type array_5bit is array(0 to 31) of std_logic_vector (4 downto 0);
end array_5bit;